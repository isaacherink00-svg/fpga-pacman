`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/20/2024 09:17:47 PM
// Design Name: 
// Module Name: maze_memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*
module maze_memory (
    input  logic [9:0]  maze_address,
    output logic [0:0]  maze_data,
    input logic clk_25MHz
);
    // Instantiate the BRAM
    maze_bram maze_bram_inst (
        .clka(clk_25MHz),
 //       .wea(1'b0),
        .addra(address),
  //      .dina(1'b0),
        .douta(maze_data)
    );
endmodule

*/